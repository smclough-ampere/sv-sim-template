module main;
  initial begin
    $display("Hello, world!");
  end
endmodule

